library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gba_bios is
   port
   (
      clk       : in std_logic;
      address   : in std_logic_vector(11 downto 0);
      data      : out std_logic_vector(31 downto 0);

      wraddress : in std_logic_vector(11 downto 0);
      wrdata    : in std_logic_vector(31 downto 0);
      wren      : in std_logic
   );
end entity;

architecture arch of gba_bios is

   type t_rom is array(0 to 4095) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"EA00000C",
      x"EA000015",
      x"EA000015",
      x"EA000013",
      x"EA000012",
      x"EA000011",
      x"EA000000",
      x"EAFFFFFF",
      x"E92D500F",
      x"E3A00301",
      x"E1A0E00F",
      x"E510F004",
      x"E8BD500F",
      x"E25EF004",
      x"E3A000DF",
      x"E129F000",
      x"E3A03301",
      x"E5C33208",
      x"EB0005F8",
      x"E3A02001",
      x"E5C32208",
      x"E59F0104",
      x"E59FE104",
      x"E12FFF10",
      x"EAFFFFFE",
      x"E92D5800",
      x"E55EC002",
      x"E28FB03C",
      x"E79BC10C",
      x"E14FB000",
      x"E92D0800",
      x"E20BB080",
      x"E38BB01F",
      x"E129F00B",
      x"E92D400C",
      x"E28FE000",
      x"E12FFF1C",
      x"E8BD400C",
      x"E3A0C0D3",
      x"E129F00C",
      x"E8BD0800",
      x"E169F00B",
      x"E8BD5800",
      x"E1B0F00E",
      x"00001804",
      x"00001524",
      x"000003D8",
      x"000003E8",
      x"00000434",
      x"000004D4",
      x"000017A8",
      x"00001798",
      x"000004E0",
      x"000004E4",
      x"0000056C",
      x"00000614",
      x"00000720",
      x"000007D8",
      x"000007E4",
      x"000008E0",
      x"00000984",
      x"00000A44",
      x"00000CDC",
      x"00000CE4",
      x"00000F18",
      x"00000FBC",
      x"000010C0",
      x"0000111C",
      x"000011AC",
      x"0000015C",
      x"0000015C",
      x"0000015C",
      x"0000015C",
      x"0000015C",
      x"0000015C",
      x"00001218",
      x"0000015C",
      x"0000015C",
      x"0000015C",
      x"00001500",
      x"00001504",
      x"0000015C",
      x"0000015C",
      x"000003CC",
      x"0000015C",
      x"0000015C",
      x"00001508",
      x"E12FFF1E",
      x"000001B8",
      x"00001804",
      x"E1A00000",
      x"E1A00000",
      x"E0832190",
      x"E1A00003",
      x"E12FFF1E",
      x"E3520000",
      x"012FFF1E",
      x"E1A03000",
      x"E0631001",
      x"E0800082",
      x"E3E0C4F1",
      x"E153000C",
      x"91D320B0",
      x"859F2010",
      x"E18120B3",
      x"E2833002",
      x"E1530000",
      x"1AFFFFF8",
      x"E12FFF1E",
      x"00001CAD",
      x"E92D4008",
      x"E59FE09C",
      x"E59FC09C",
      x"E1A0200E",
      x"E3A03405",
      x"E3E004F1",
      x"E1520000",
      x"908E1003",
      x"928114FB",
      x"91D110B0",
      x"859F1080",
      x"E0C310B2",
      x"E153000C",
      x"E2822002",
      x"1AFFFFF6",
      x"E59F0070",
      x"E3A01406",
      x"E3A02000",
      x"EB000255",
      x"E59F1064",
      x"E3A02000",
      x"E59F0060",
      x"EB000251",
      x"E3A03301",
      x"E3A02C1E",
      x"E1C320B8",
      x"E3A02C01",
      x"E5832000",
      x"E3A01077",
      x"E1D320B6",
      x"E352009F",
      x"8AFFFFFC",
      x"E1D320B6",
      x"E352009F",
      x"9AFFFFFC",
      x"E3510000",
      x"E2411001",
      x"1AFFFFF6",
      x"E3A000FF",
      x"EB0004B2",
      x"E8BD4008",
      x"E12FFF1E",
      x"00001888",
      x"05000040",
      x"00001CAD",
      x"00001A98",
      x"0600F000",
      x"000018A8",
      x"E3500000",
      x"B3E03000",
      x"A3A03000",
      x"E0830000",
      x"E0200003",
      x"E12FFF1E",
      x"E3700107",
      x"82800103",
      x"83A02205",
      x"93A02201",
      x"83A03801",
      x"93A03000",
      x"E1500002",
      x"23833902",
      x"20620000",
      x"E2832A02",
      x"E1A02682",
      x"E1500002",
      x"23833901",
      x"20620000",
      x"E2832A01",
      x"E1A02602",
      x"E1500002",
      x"23833A02",
      x"20620000",
      x"E2832B02",
      x"E1A02582",
      x"E1500002",
      x"23833A01",
      x"20620000",
      x"E2832B01",
      x"E1A02502",
      x"E1500002",
      x"23833B02",
      x"20620000",
      x"E2832C02",
      x"E1A02482",
      x"E1500002",
      x"23833B01",
      x"20620000",
      x"E2832C01",
      x"E1A02402",
      x"E1500002",
      x"23833C02",
      x"20620000",
      x"E2832080",
      x"E1A02382",
      x"E1500002",
      x"23833C01",
      x"20620000",
      x"E2832040",
      x"E1A02302",
      x"E1500002",
      x"23833080",
      x"20620000",
      x"E2832020",
      x"E1A02282",
      x"E1500002",
      x"23833040",
      x"20620000",
      x"E2832010",
      x"E1A02202",
      x"E1500002",
      x"23833020",
      x"20620000",
      x"E2832008",
      x"E1A02182",
      x"E1500002",
      x"23833010",
      x"20620000",
      x"E2832004",
      x"E1A02102",
      x"E1500002",
      x"23833008",
      x"20620000",
      x"E2832002",
      x"E1A02082",
      x"E1500002",
      x"23833004",
      x"20620000",
      x"E2832001",
      x"E1500002",
      x"23833002",
      x"E1A000A3",
      x"E12FFF1E",
      x"E3A03301",
      x"E5C30301",
      x"E12FFF1E",
      x"E3A02000",
      x"E3A03301",
      x"E5C32301",
      x"E12FFF1E",
      x"E3E0207F",
      x"E3A03301",
      x"E5C32301",
      x"E12FFF1E",
      x"E3A01000",
      x"E3A03F82",
      x"E3A02301",
      x"E18210B3",
      x"E3E0233F",
      x"E15230B7",
      x"E0130000",
      x"10203003",
      x"114230B7",
      x"E3A01001",
      x"E3A03F82",
      x"E3A02301",
      x"E20000FF",
      x"E18210B3",
      x"E12FFF1E",
      x"E3500000",
      x"01A01801",
      x"E92D00F0",
      x"01A00821",
      x"0A00000E",
      x"E3A00000",
      x"E3A03F82",
      x"E3A02301",
      x"E18200B3",
      x"E3E0233F",
      x"E15230B7",
      x"E1A01801",
      x"E1A00821",
      x"E0101003",
      x"10213003",
      x"114230B7",
      x"E3A01001",
      x"E3A03F82",
      x"E3A02301",
      x"E18210B3",
      x"E3A05000",
      x"E3A02301",
      x"E3A0CF82",
      x"E1A07005",
      x"E3E0433F",
      x"E3A06001",
      x"E5C25301",
      x"E18270BC",
      x"E15430B7",
      x"E0101003",
      x"E0213003",
      x"0A000005",
      x"E31100FF",
      x"E14430B7",
      x"E18260BC",
      x"0AFFFFF5",
      x"E8BD00F0",
      x"E12FFF1E",
      x"E18260BC",
      x"EAFFFFF1",
      x"E3A00001",
      x"E1A01000",
      x"EAFFFFD4",
      x"EAFFFF6A",
      x"E0030090",
      x"E1A03743",
      x"E2633000",
      x"E0832083",
      x"E0622182",
      x"E0832182",
      x"E1A02742",
      x"E2822E39",
      x"E0020293",
      x"E1A02742",
      x"E2822E91",
      x"E282200C",
      x"E0020293",
      x"E1A02742",
      x"E2822EFB",
      x"E2822006",
      x"E0020293",
      x"E1A02742",
      x"E2822D5A",
      x"E282202A",
      x"E0020293",
      x"E1A02742",
      x"E2822D82",
      x"E0223293",
      x"E1A02742",
      x"E2822DD9",
      x"E2822011",
      x"E0030392",
      x"E1A03743",
      x"E2833CA2",
      x"E28330F9",
      x"E0000093",
      x"E1A00840",
      x"E12FFF1E",
      x"E92D4038",
      x"E2515000",
      x"E1A04000",
      x"01A04840",
      x"02040902",
      x"0A000010",
      x"E3540000",
      x"0A000010",
      x"E0242FC4",
      x"E0422FC4",
      x"E0253FC5",
      x"E0433FC5",
      x"E1520003",
      x"CA000011",
      x"0A00000D",
      x"E1A01005",
      x"E1A00704",
      x"EB00047C",
      x"EBFFFFCA",
      x"E1A04845",
      x"E2044902",
      x"E2844901",
      x"E0600004",
      x"E8BD4038",
      x"E12FFF1E",
      x"E1A00845",
      x"E2000902",
      x"E2800901",
      x"EAFFFFF9",
      x"E3540000",
      x"B3550000",
      x"BAFFFFEE",
      x"E1A00705",
      x"E1A01004",
      x"EB00046B",
      x"EBFFFFB9",
      x"E3540000",
      x"A1A057A5",
      x"A2055801",
      x"B2800902",
      x"A0800005",
      x"EAFFFFEC",
      x"E310040E",
      x"E52D4004",
      x"0A000018",
      x"E1A03582",
      x"E1A034A3",
      x"E3C3360E",
      x"E0833000",
      x"E313040E",
      x"0A000012",
      x"E3C234FF",
      x"E3120301",
      x"E3C3360E",
      x"1A000010",
      x"E3120401",
      x"1A00001E",
      x"E3530000",
      x"0A00000A",
      x"E1A02000",
      x"E0803083",
      x"E0601001",
      x"E3E044F1",
      x"E1520004",
      x"91D2C0B0",
      x"859FC0A0",
      x"E181C0B2",
      x"E2822002",
      x"E1520003",
      x"1AFFFFF8",
      x"E8BD0010",
      x"E12FFF1E",
      x"E3120401",
      x"E3C11003",
      x"E3C02003",
      x"1A000015",
      x"E3530000",
      x"10621001",
      x"13E0C4F1",
      x"0AFFFFF5",
      x"E152000C",
      x"95920000",
      x"859F0060",
      x"E2533001",
      x"E7810002",
      x"E2822004",
      x"1AFFFFF8",
      x"EAFFFFED",
      x"E350040F",
      x"31D020B0",
      x"259F203C",
      x"E3530000",
      x"0AFFFFE8",
      x"E0813083",
      x"E0C120B2",
      x"E1510003",
      x"1AFFFFFC",
      x"EAFFFFE3",
      x"E352040F",
      x"35922000",
      x"259F2018",
      x"E3530000",
      x"0AFFFFDE",
      x"E2533001",
      x"E4812004",
      x"1AFFFFFC",
      x"EAFFFFDA",
      x"00001CAD",
      x"1CAD1CAD",
      x"E310040E",
      x"E52D4004",
      x"0A000017",
      x"E1A03582",
      x"E1A034A3",
      x"E3C3360E",
      x"E0833000",
      x"E313040E",
      x"0A000011",
      x"E3C244FF",
      x"E3120401",
      x"E3C03003",
      x"E3C11003",
      x"E3C4460E",
      x"0A00000D",
      x"E353040F",
      x"35932000",
      x"259F2068",
      x"E3540000",
      x"0A000006",
      x"E2813020",
      x"E4812004",
      x"E1510003",
      x"1AFFFFFC",
      x"E2444008",
      x"E3540000",
      x"CAFFFFF8",
      x"E8BD0010",
      x"E12FFF1E",
      x"E3540000",
      x"10631001",
      x"13E0C4F1",
      x"0AFFFFF9",
      x"E2830020",
      x"E153000C",
      x"95932000",
      x"859F201C",
      x"E7812003",
      x"E2833004",
      x"E1530000",
      x"1AFFFFF8",
      x"E2444008",
      x"E3540000",
      x"CAFFFFF4",
      x"EAFFFFED",
      x"BAFFFFFB",
      x"E59F0000",
      x"E12FFF1E",
      x"BAAE187F",
      x"E3520000",
      x"E92D0FF0",
      x"E2422001",
      x"0A000037",
      x"E2800014",
      x"E2811010",
      x"E150C0B4",
      x"E1A0C42C",
      x"E28C3040",
      x"E59F40CC",
      x"E20330FF",
      x"E1A03083",
      x"E15060F8",
      x"E19430F3",
      x"E0040693",
      x"E59F70B4",
      x"E1A0C08C",
      x"E15080F6",
      x"E19750FC",
      x"E00C0895",
      x"E15070BC",
      x"E1A04744",
      x"E0030398",
      x"E0050596",
      x"E1A07807",
      x"E1A0A804",
      x"E1A07847",
      x"E1A0A84A",
      x"E00A0A97",
      x"E1A0C74C",
      x"E15060BA",
      x"E1A0B80C",
      x"E1A03743",
      x"E1A0B84B",
      x"E1A05745",
      x"E00B0B97",
      x"E1A06806",
      x"E5107014",
      x"E1A09803",
      x"E1A06846",
      x"E1A08805",
      x"E1A09849",
      x"E06AA007",
      x"E0090996",
      x"E1A08848",
      x"E026A698",
      x"E5107010",
      x"E2422001",
      x"E06B7007",
      x"E2655000",
      x"E0697007",
      x"E3720001",
      x"E14141B0",
      x"E14150BE",
      x"E141C0BC",
      x"E14130BA",
      x"E90100C0",
      x"E2800014",
      x"E2811010",
      x"1AFFFFC9",
      x"E8BD0FF0",
      x"E12FFF1E",
      x"00002150",
      x"E3520000",
      x"E92D07F0",
      x"E2422001",
      x"0A000021",
      x"E1A07083",
      x"E59FA084",
      x"E0878083",
      x"E2800008",
      x"E0813003",
      x"E150C0B4",
      x"E1A0C42C",
      x"E28C4040",
      x"E20440FF",
      x"E1A0C08C",
      x"E15060F8",
      x"E19A50FC",
      x"E1A0C084",
      x"E19AC0FC",
      x"E15040F6",
      x"E0090596",
      x"E006069C",
      x"E0050594",
      x"E00C0C94",
      x"E1A09749",
      x"E2422001",
      x"E1A06746",
      x"E2699000",
      x"E1A05745",
      x"E1A0C74C",
      x"E3720001",
      x"E1C160B0",
      x"E2800008",
      x"E1C390B0",
      x"E18150B7",
      x"E183C0B7",
      x"E0811008",
      x"E0833008",
      x"1AFFFFE2",
      x"E8BD07F0",
      x"E12FFF1E",
      x"00002150",
      x"E92D0FF0",
      x"E310040E",
      x"E24DD008",
      x"E1D2C0B0",
      x"0A000027",
      x"E08CC000",
      x"E31C040E",
      x"0A000024",
      x"E5D27002",
      x"E3A050FF",
      x"E2673008",
      x"E1A05355",
      x"E5923004",
      x"E3A06000",
      x"E5D2B003",
      x"E150000C",
      x"E1A02FA3",
      x"E3C33102",
      x"E58D2000",
      x"E58D3004",
      x"E1A0A006",
      x"0A000016",
      x"E4D04001",
      x"E1A02005",
      x"E3A03000",
      x"E59D8000",
      x"E0029004",
      x"E3590000",
      x"13888001",
      x"E3580000",
      x"E1A08339",
      x"159D9004",
      x"10888009",
      x"E18AA618",
      x"E086600B",
      x"E356001F",
      x"C3A06000",
      x"E0833007",
      x"C481A004",
      x"C1A0A006",
      x"E3530007",
      x"E1A02712",
      x"DAFFFFED",
      x"E150000C",
      x"1AFFFFE8",
      x"E28DD008",
      x"E8BD0FF0",
      x"E12FFF1E",
      x"E4902004",
      x"E310040E",
      x"E92D01F0",
      x"0A00001C",
      x"E1A02422",
      x"E3C234FF",
      x"E3C3360E",
      x"E0833000",
      x"E313040E",
      x"0A000016",
      x"E3520000",
      x"0A000014",
      x"E5D04000",
      x"E3540000",
      x"E280C001",
      x"0A000012",
      x"E3A08008",
      x"E3140080",
      x"1A00001A",
      x"E5DC3000",
      x"E2522001",
      x"E2810001",
      x"E28CC001",
      x"E5C13000",
      x"0A000007",
      x"E1A01000",
      x"E1A04084",
      x"E2588001",
      x"E20440FF",
      x"1AFFFFF2",
      x"E3520000",
      x"E1A0000C",
      x"CAFFFFEA",
      x"E8BD01F0",
      x"E12FFF1E",
      x"E2804009",
      x"E1A0000C",
      x"E4D03001",
      x"E2522001",
      x"E4C13001",
      x"0AFFFFF7",
      x"E1500004",
      x"1AFFFFF9",
      x"E3520000",
      x"CAFFFFDE",
      x"EAFFFFF2",
      x"E5DC0000",
      x"E5DC3001",
      x"E1833400",
      x"E1A03803",
      x"E1A07E23",
      x"E2416001",
      x"E1A03203",
      x"E2420001",
      x"E0466A23",
      x"E2877003",
      x"E1A05000",
      x"E3A03000",
      x"EA000000",
      x"E2400001",
      x"E7D32006",
      x"E1530005",
      x"E4C12001",
      x"E2833001",
      x"E1A02000",
      x"0AFFFFDE",
      x"E1570003",
      x"CAFFFFF6",
      x"E28CC002",
      x"EAFFFFD3",
      x"E92D0FF0",
      x"E4905004",
      x"E3520000",
      x"01A05425",
      x"0A000007",
      x"E310040E",
      x"0A000024",
      x"E1A05425",
      x"E3C534FF",
      x"E3C3360E",
      x"E0833000",
      x"E313040E",
      x"0A00001E",
      x"E3550000",
      x"0A00001C",
      x"E3A03000",
      x"E1A0C003",
      x"E1A04003",
      x"E5D07000",
      x"E3570000",
      x"E2806001",
      x"0A000017",
      x"E3A0B008",
      x"E3170080",
      x"1A000026",
      x"E5D62000",
      x"E1833C12",
      x"E3540001",
      x"00C130B2",
      x"03A03000",
      x"128CC008",
      x"13A04001",
      x"01A0C003",
      x"01A04003",
      x"E2555001",
      x"E2866001",
      x"0A000006",
      x"E1A07087",
      x"E25BB001",
      x"E20770FF",
      x"1AFFFFED",
      x"E3550000",
      x"E1A00006",
      x"CAFFFFE5",
      x"E8BD0FF0",
      x"E12FFF1E",
      x"E2807009",
      x"E1A00006",
      x"E4D02001",
      x"E1833C12",
      x"E3540001",
      x"00C130B2",
      x"03A03000",
      x"128CC008",
      x"13A04001",
      x"01A0C003",
      x"01A04003",
      x"E2555001",
      x"0AFFFFF0",
      x"E1500007",
      x"1AFFFFF2",
      x"E3550000",
      x"CAFFFFD2",
      x"EAFFFFEB",
      x"E5D60000",
      x"E5D62001",
      x"E1822400",
      x"E1A02802",
      x"E241A001",
      x"E1A09E22",
      x"E08AA004",
      x"E1A02202",
      x"E2450001",
      x"E04AAA22",
      x"E2899003",
      x"E1A08000",
      x"E3A02000",
      x"EA000000",
      x"E2400001",
      x"E7D2500A",
      x"E1833C15",
      x"E3540001",
      x"00C130B2",
      x"03A03000",
      x"128CC008",
      x"13A04001",
      x"01A0C003",
      x"01A04003",
      x"E1520008",
      x"E1A05000",
      x"E2822001",
      x"0AFFFFCF",
      x"E1590002",
      x"CAFFFFEF",
      x"E2866002",
      x"EAFFFFC4",
      x"E3A02001",
      x"EAFFFF9D",
      x"E92D0FF0",
      x"E1A03000",
      x"E4934004",
      x"E24DD010",
      x"E313040E",
      x"E58D1000",
      x"0A000033",
      x"E1A02424",
      x"E3C214FF",
      x"E3C1160E",
      x"E0813003",
      x"E313040E",
      x"0A00002D",
      x"E5D0C004",
      x"E2806005",
      x"E28CC001",
      x"E204400F",
      x"E086C08C",
      x"E3540008",
      x"E51C3001",
      x"E5D07005",
      x"E28CC003",
      x"0A000048",
      x"E3520000",
      x"DA000021",
      x"E3A08000",
      x"E58D800C",
      x"E58D8004",
      x"E58D8008",
      x"E1A05007",
      x"E1A09008",
      x"E3A01102",
      x"E3A04001",
      x"E1110003",
      x"11A05325",
      x"1084B000",
      x"1205A001",
      x"01A0A3A5",
      x"15DB5006",
      x"07D45006",
      x"E35A0000",
      x"0A000005",
      x"E3590000",
      x"1A000011",
      x"E1888005",
      x"E3A09004",
      x"E1A05007",
      x"E3A04000",
      x"E1B010A1",
      x"049C3004",
      x"03A01102",
      x"E3520000",
      x"DA000005",
      x"E3540000",
      x"0AFFFFE8",
      x"E205A03F",
      x"E28AA001",
      x"E084408A",
      x"EAFFFFE5",
      x"E28DD010",
      x"E8BD0FF0",
      x"E12FFF1E",
      x"E2899004",
      x"E3590008",
      x"E1888205",
      x"13A04000",
      x"11A05007",
      x"1AFFFFEB",
      x"E59D5004",
      x"E2855001",
      x"E59D400C",
      x"E58D5004",
      x"E3550004",
      x"E59D5008",
      x"E1844518",
      x"E3A08000",
      x"E58D400C",
      x"0A000005",
      x"E2855008",
      x"E58D5008",
      x"E1A09008",
      x"E1A05007",
      x"E1A04008",
      x"EAFFFFDB",
      x"E59D5000",
      x"E59D400C",
      x"E4854004",
      x"E2422004",
      x"E58D5000",
      x"E1A09008",
      x"E1A05007",
      x"E58D800C",
      x"E58D8004",
      x"E58D8008",
      x"E1A04008",
      x"EAFFFFCF",
      x"E3520000",
      x"DAFFFFD8",
      x"E3A0A000",
      x"E1A05007",
      x"E3A01102",
      x"E1A0B00A",
      x"E1A0900A",
      x"E3A04001",
      x"E1130001",
      x"11A08325",
      x"01A083A5",
      x"10845000",
      x"12088001",
      x"15D55006",
      x"07D45006",
      x"E3580000",
      x"0A000006",
      x"E2899001",
      x"E3590004",
      x"E18AAB15",
      x"0A00000D",
      x"E28BB008",
      x"E1A05007",
      x"E3A04000",
      x"E1B010A1",
      x"049C3004",
      x"03A01102",
      x"E3520000",
      x"DAFFFFBD",
      x"E3540000",
      x"0AFFFFE7",
      x"E205803F",
      x"E2888001",
      x"E0844088",
      x"EAFFFFE4",
      x"E59D4000",
      x"E484A004",
      x"E3A0A000",
      x"E58D4000",
      x"E2422004",
      x"E1A05007",
      x"E1A0900A",
      x"E1A0B00A",
      x"E1A0400A",
      x"EAFFFFEA",
      x"E4902004",
      x"E310040E",
      x"E92D0030",
      x"0A000017",
      x"E1A02422",
      x"E3C234FF",
      x"E3C3360E",
      x"E0833000",
      x"E313040E",
      x"0A000011",
      x"E3520000",
      x"0A00000F",
      x"E5D04000",
      x"E3140080",
      x"E280C001",
      x"E204407F",
      x"01A03001",
      x"1A00000B",
      x"E4DC0001",
      x"E4C30001",
      x"E2522001",
      x"E0610003",
      x"0A000004",
      x"E1540000",
      x"AAFFFFF8",
      x"E1A01003",
      x"E1A0000C",
      x"EAFFFFEF",
      x"E8BD0030",
      x"E12FFF1E",
      x"E5D05001",
      x"E2844003",
      x"E1A03001",
      x"E4C35001",
      x"E2522001",
      x"E061C003",
      x"0AFFFFF6",
      x"E154000C",
      x"CAFFFFF9",
      x"E280C002",
      x"EAFFFFEF",
      x"E92D05F0",
      x"E2806004",
      x"E316040E",
      x"E3C00003",
      x"E5900000",
      x"0A000021",
      x"E1A00420",
      x"E3C034FF",
      x"E3C3360E",
      x"E0833006",
      x"E313040E",
      x"0A00001B",
      x"E3500000",
      x"0A000019",
      x"E3A03000",
      x"E1A02003",
      x"E1A04003",
      x"E5D67000",
      x"E3170080",
      x"E2865001",
      x"E207707F",
      x"03A0C000",
      x"1A000012",
      x"E4D56001",
      x"E1833216",
      x"E3540001",
      x"00C130B2",
      x"03A03000",
      x"12822008",
      x"13A04001",
      x"01A02003",
      x"01A04003",
      x"E2500001",
      x"E28CC001",
      x"0A000004",
      x"E157000C",
      x"AAFFFFF1",
      x"E1A06005",
      x"E3500000",
      x"CAFFFFE8",
      x"E8BD05F0",
      x"E12FFF1E",
      x"E2405001",
      x"E5D6A001",
      x"E2877003",
      x"E1A08005",
      x"E3A0C000",
      x"EA000000",
      x"E2455001",
      x"E183321A",
      x"E3540001",
      x"00C130B2",
      x"03A03000",
      x"12822008",
      x"13A04001",
      x"01A02003",
      x"01A04003",
      x"E15C0008",
      x"E1A00005",
      x"E28CC001",
      x"0AFFFFEA",
      x"E157000C",
      x"CAFFFFF0",
      x"E2866002",
      x"EAFFFFE4",
      x"E1A02000",
      x"E492C004",
      x"E312040E",
      x"012FFF1E",
      x"E1A0C42C",
      x"E3CC34FF",
      x"E3C3360E",
      x"E0833002",
      x"E313040E",
      x"012FFF1E",
      x"E5D03004",
      x"E35C0001",
      x"E2800005",
      x"E5C13000",
      x"D12FFF1E",
      x"E082C00C",
      x"E4D02001",
      x"E0833002",
      x"E20330FF",
      x"E150000C",
      x"E5E13001",
      x"1AFFFFF9",
      x"E12FFF1E",
      x"E1A03000",
      x"E92D0070",
      x"E4936004",
      x"E313040E",
      x"0A00001C",
      x"E1A06426",
      x"E3C624FF",
      x"E3C2260E",
      x"E0823003",
      x"E313040E",
      x"0A000016",
      x"E5D03004",
      x"E3560001",
      x"E2800005",
      x"E1A0C003",
      x"DA000011",
      x"E3A04001",
      x"E3A02008",
      x"E4D05001",
      x"E0833005",
      x"E20330FF",
      x"E18CC213",
      x"E3540001",
      x"E1A0C80C",
      x"03A04000",
      x"E1A0C82C",
      x"02466002",
      x"00C1C0B2",
      x"12822008",
      x"13A04001",
      x"01A02004",
      x"01A0C004",
      x"E3560001",
      x"CAFFFFEF",
      x"E8BD0070",
      x"E12FFF1E",
      x"E1A03000",
      x"E493C004",
      x"E313040E",
      x"012FFF1E",
      x"E1A0C42C",
      x"E3CC24FF",
      x"E3C2260E",
      x"E0823003",
      x"E313040E",
      x"012FFF1E",
      x"E1D030B4",
      x"E35C0003",
      x"E2802006",
      x"E1C130B0",
      x"D12FFF1E",
      x"E24CC004",
      x"E2800008",
      x"E3CCC001",
      x"E080C00C",
      x"E0D200B2",
      x"E0833000",
      x"E1A03803",
      x"E1A03823",
      x"E152000C",
      x"E1E130B2",
      x"1AFFFFF8",
      x"E12FFF1E",
      x"E35100B2",
      x"E92D4038",
      x"E59F3064",
      x"83A010B2",
      x"E1A05000",
      x"92810001",
      x"E0831001",
      x"E5D1C200",
      x"E20C100F",
      x"E0831101",
      x"E59142B4",
      x"E1A0C22C",
      x"E1A04C34",
      x"83A000B3",
      x"E0831000",
      x"E5D1C200",
      x"E20C100F",
      x"E0833101",
      x"E59302B4",
      x"83A024FF",
      x"E1A0C22C",
      x"E1A01002",
      x"E0640C30",
      x"EBFFFBBD",
      x"E5951004",
      x"E0840000",
      x"EBFFFBBA",
      x"E8BD4038",
      x"E12FFF1E",
      x"00002150",
      x"E59F325C",
      x"E92D47F0",
      x"E5934FF0",
      x"E59F3254",
      x"E5942000",
      x"E1520003",
      x"0A000001",
      x"E8BD47F0",
      x"E12FFF1E",
      x"E5943020",
      x"E59F223C",
      x"E3530000",
      x"E5842000",
      x"15940024",
      x"11A0E00F",
      x"112FFF13",
      x"E5943028",
      x"E3530000",
      x"15940024",
      x"11A0E00F",
      x"112FFF13",
      x"E5D42004",
      x"E3520000",
      x"E2843E35",
      x"E5940010",
      x"0A000076",
      x"E5D4100B",
      x"E2811001",
      x"E0621001",
      x"E20110FF",
      x"E0213190",
      x"E5D46005",
      x"E3560000",
      x"02812E63",
      x"01A08001",
      x"0A000018",
      x"E3520002",
      x"0A000000",
      x"E0813000",
      x"E2807001",
      x"E5D1C000",
      x"E2812E63",
      x"E1A08001",
      x"E0877003",
      x"E1D290D0",
      x"E2835E63",
      x"E1D5A0D0",
      x"E1A0CC0C",
      x"E0D350D1",
      x"E089CC4C",
      x"E08CC00A",
      x"E08CC005",
      x"E00C0C96",
      x"E1A0C4CC",
      x"E31C0080",
      x"128CC001",
      x"E20CC0FF",
      x"E1530007",
      x"E5C2C000",
      x"E5C1C000",
      x"1AFFFFEE",
      x"E1B031A0",
      x"1A00004D",
      x"E2810E63",
      x"E5883000",
      x"E281C004",
      x"E5823000",
      x"E2802004",
      x"E3A03000",
      x"E58C3000",
      x"E28C1008",
      x"E5823000",
      x"E1A00003",
      x"E58C3004",
      x"E5823004",
      x"E2822008",
      x"E2811010",
      x"E2822010",
      x"E3A03000",
      x"E2400001",
      x"E3700001",
      x"E5013010",
      x"E5023010",
      x"E501300C",
      x"E502300C",
      x"E5013008",
      x"E5023008",
      x"E5013004",
      x"E5023004",
      x"E2811010",
      x"E2822010",
      x"1AFFFFF2",
      x"E5D47006",
      x"E2846090",
      x"E1A03006",
      x"E1A02007",
      x"E3A08003",
      x"E3A05000",
      x"E5531040",
      x"E31100C7",
      x"E513001C",
      x"0A00001E",
      x"E3110080",
      x"1A00001C",
      x"E3110040",
      x"E280C010",
      x"0A000019",
      x"E5438040",
      x"E503C018",
      x"E590000C",
      x"E5030028",
      x"E553003C",
      x"E31100C0",
      x"03A0C003",
      x"13A0C013",
      x"E35000FF",
      x"E1A0100C",
      x"024C1001",
      x"020110FF",
      x"E5435037",
      x"E543C040",
      x"E5035024",
      x"05431040",
      x"E5430037",
      x"E5D40007",
      x"E0211190",
      x"E553003E",
      x"E1A01201",
      x"E0010190",
      x"E1A01421",
      x"E20110FF",
      x"E5431036",
      x"E5431035",
      x"E2422001",
      x"E20220FF",
      x"E35200FF",
      x"E2833040",
      x"1AFFFFD7",
      x"E59F3038",
      x"E7863307",
      x"EAFFFF79",
      x"E1B00220",
      x"1AFFFFBC",
      x"E1A0C001",
      x"EAFFFFB2",
      x"E5D46005",
      x"E3560000",
      x"01A08003",
      x"02842D26",
      x"01A01003",
      x"0AFFFFA5",
      x"E1A01003",
      x"EAFFFF8C",
      x"03007000",
      x"68736D53",
      x"68736D54",
      x"E12FFF1E",
      x"E12FFF1E",
      x"E59F2010",
      x"E2803090",
      x"E4802004",
      x"E1500003",
      x"1AFFFFFC",
      x"E12FFF1E",
      x"0000015C",
      x"E92D4010",
      x"E3A03000",
      x"E24DD008",
      x"E58D3004",
      x"E3A02080",
      x"E3A03301",
      x"E2504000",
      x"E1C320B0",
      x"0A000064",
      x"E3140001",
      x"1A00006C",
      x"E3140002",
      x"1A000070",
      x"E3140004",
      x"1A000074",
      x"E3140008",
      x"1A000078",
      x"E3140010",
      x"1A00005D",
      x"E3140080",
      x"0A000020",
      x"E59F31E8",
      x"E59F11E8",
      x"E3A02000",
      x"E1E320B2",
      x"E1530001",
      x"1AFFFFFC",
      x"E59F11D8",
      x"E3A03381",
      x"E3A02000",
      x"E1E320B2",
      x"E1530001",
      x"1AFFFFFC",
      x"E59F31C4",
      x"E59F11C4",
      x"E3A02000",
      x"E1E320B2",
      x"E1530001",
      x"1AFFFFFC",
      x"E59F31B4",
      x"E59F11B4",
      x"E3A02000",
      x"E1E320B2",
      x"E1530001",
      x"1AFFFFFC",
      x"E3A03301",
      x"E3A02C01",
      x"E3A01E13",
      x"E3A00000",
      x"E18300B1",
      x"E1C322B0",
      x"E1C323B0",
      x"E1C322B6",
      x"E1C323B6",
      x"E3140020",
      x"0A000022",
      x"E3A03301",
      x"E3A02000",
      x"E3A01E11",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A01F45",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A01F46",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A01F47",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A00902",
      x"E3A01F4D",
      x"E18300B1",
      x"E3A01D05",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A01F51",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A01F52",
      x"E18320B1",
      x"E2811002",
      x"E18320B1",
      x"E3A01F53",
      x"E18320B1",
      x"E3140040",
      x"0A000010",
      x"E3A03301",
      x"E1D318B8",
      x"E59F00DC",
      x"E3A02000",
      x"E3C11B3F",
      x"E5830080",
      x"E1C318B8",
      x"E5C32070",
      x"E1C329B0",
      x"E1C329B2",
      x"E1C329B4",
      x"E1C329B6",
      x"E1C329B8",
      x"E1C329BA",
      x"E1C329BC",
      x"E1C329BE",
      x"E5C32084",
      x"E28DD008",
      x"E8BD4010",
      x"E12FFF1E",
      x"E28D0004",
      x"E3A01407",
      x"E59F2090",
      x"EBFFFC09",
      x"E3140080",
      x"0AFFFFBE",
      x"EAFFFF9C",
      x"E28D0004",
      x"E3A01402",
      x"E59F2078",
      x"EBFFFC02",
      x"E3140002",
      x"0AFFFF8E",
      x"E28D0004",
      x"E3A01403",
      x"E59F2064",
      x"EBFFFBFC",
      x"E3140004",
      x"0AFFFF8A",
      x"E28D0004",
      x"E3A01405",
      x"E59F2044",
      x"EBFFFBF6",
      x"E3140008",
      x"0AFFFF86",
      x"E28D0004",
      x"E3A01406",
      x"E59F2038",
      x"EBFFFBF0",
      x"E3140010",
      x"0AFFFF82",
      x"EAFFFFDF",
      x"040001FE",
      x"0400021E",
      x"04000020",
      x"0400001E",
      x"0400005E",
      x"040000AE",
      x"040000DE",
      x"880E0000",
      x"01000100",
      x"01010000",
      x"01001F80",
      x"01006000",
      x"E1A03000",
      x"E1A00001",
      x"E1A01003",
      x"EAFFFFFF",
      x"E210C102",
      x"42600000",
      x"E2113102",
      x"42611000",
      x"E02CC003",
      x"E3A02000",
      x"E3A03001",
      x"E1510000",
      x"91A01081",
      x"91A03083",
      x"9AFFFFFB",
      x"E1500001",
      x"20400001",
      x"21822003",
      x"E1B030A3",
      x"31A010A1",
      x"3AFFFFF9",
      x"E1A01000",
      x"E1A03002",
      x"E1A00002",
      x"E31C0102",
      x"42600000",
      x"E12FFF1E",
      x"E3A03301",
      x"E5532006",
      x"EB000007",
      x"E3520000",
      x"E9131FFF",
      x"13A0E402",
      x"03A0E302",
      x"E3A0001F",
      x"E129F000",
      x"E3A00000",
      x"E12FFF1E",
      x"E3A000D3",
      x"E129F000",
      x"E59FD044",
      x"E3A0E000",
      x"E169F00E",
      x"E3A000D2",
      x"E129F000",
      x"E59FD02C",
      x"E3A0E000",
      x"E169F00E",
      x"E3A0005F",
      x"E129F000",
      x"E59FD014",
      x"E3B00000",
      x"E2501C02",
      x"E7830001",
      x"E2911004",
      x"BAFFFFFC",
      x"E12FFF1E",
      x"03007F00",
      x"03007FA0",
      x"03007FE0",
      x"04210000",
      x"0C630842",
      x"18C61084",
      x"21081CE7",
      x"2D6B294A",
      x"63184631",
      x"77BD6F7B",
      x"7FFF7BDE",
      x"00080010",
      x"F000003F",
      x"F001F001",
      x"F001F001",
      x"FF01F001",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"F001F0FF",
      x"F001F001",
      x"F001F001",
      x"7001F001",
      x"00011D07",
      x"F001F002",
      x"030B4001",
      x"040140A0",
      x"06000500",
      x"01F00700",
      x"4001F0C1",
      x"0900080B",
      x"84400A00",
      x"0C000B00",
      x"0E000D00",
      x"000F0600",
      x"F0110010",
      x"1205A098",
      x"00130002",
      x"00150014",
      x"00081619",
      x"20180017",
      x"1A001921",
      x"1B290080",
      x"1D001C00",
      x"00001E00",
      x"0020001F",
      x"00220021",
      x"24002300",
      x"26002500",
      x"00270000",
      x"00290028",
      x"2B00002A",
      x"2D002C00",
      x"00002E00",
      x"0030002F",
      x"88320031",
      x"00335B00",
      x"35612034",
      x"20803600",
      x"3800373F",
      x"3A003900",
      x"003B0000",
      x"003D003C",
      x"3F00003E",
      x"41004000",
      x"00004200",
      x"00440043",
      x"00460045",
      x"48004700",
      x"4A004900",
      x"004B0008",
      x"4D99204C",
      x"20804E00",
      x"50004FA1",
      x"52005100",
      x"00530000",
      x"00550054",
      x"57000056",
      x"59005800",
      x"00005A00",
      x"005C005B",
      x"005E005D",
      x"60005F00",
      x"62006100",
      x"00630000",
      x"00650064",
      x"67000866",
      x"D9006800",
      x"206A0069",
      x"E1406B00",
      x"006D006C",
      x"6F00386E",
      x"01F001F0",
      x"00700B40",
      x"72002071",
      x"00731F81",
      x"E3750074",
      x"01F001F0",
      x"00760B40",
      x"F05DF177",
      x"01F0FF01",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"F0FF01F0",
      x"F001F001",
      x"F001F001",
      x"F001F001",
      x"FF01F001",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"F001F0FF",
      x"F001F001",
      x"F001F001",
      x"F001F001",
      x"01F0FF01",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"F0FF01F0",
      x"F001F001",
      x"F001F001",
      x"F001F001",
      x"FF01F001",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"01F001F0",
      x"F001F0FE",
      x"F001F001",
      x"F001F001",
      x"00016001",
      x"000F0010",
      x"F000003C",
      x"F001F001",
      x"410D1001",
      x"88883376",
      x"077015F0",
      x"1FF08888",
      x"78101FA0",
      x"15F00247",
      x"00009200",
      x"00DA2000",
      x"00FFA300",
      x"FFEA2020",
      x"00951F00",
      x"00EDB940",
      x"FFFEB910",
      x"FFFFFEB7",
      x"FFFFFD14",
      x"00EF0110",
      x"06FFAB06",
      x"BA14ADFF",
      x"901030ED",
      x"AB0CCD05",
      x"40275699",
      x"FF1DF058",
      x"555508FF",
      x"77505555",
      x"C0BDEFFF",
      x"23B04700",
      x"EDCA9995",
      x"10280000",
      x"179B10A5",
      x"5ACEA000",
      x"FF000901",
      x"4B004ACF",
      x"7E0029CE",
      x"7F10AE56",
      x"938700EB",
      x"BFD00400",
      x"D000A703",
      x"CFD4005B",
      x"107B0005",
      x"A801F008",
      x"00300E10",
      x"17007013",
      x"85A200B0",
      x"FFD94300",
      x"D80060FF",
      x"80DB00B1",
      x"FBAE0A00",
      x"FE3BFFFF",
      x"04DF00FF",
      x"00AFFFFF",
      x"0401BDFF",
      x"003AFF00",
      x"44008D00",
      x"48F01862",
      x"000001F0",
      x"F01200D0",
      x"A00380C2",
      x"CDDDDD21",
      x"1A420105",
      x"8E4601AE",
      x"F0BF4A01",
      x"D0CBB03E",
      x"DD01DB02",
      x"FFFC0BDD",
      x"03500CFF",
      x"5022F0D6",
      x"63015009",
      x"501FE1F0",
      x"45755509",
      x"7DF09B01",
      x"01400680",
      x"3FF0A0A3",
      x"013F60C0",
      x"0004DF93",
      x"09FDA200",
      x"D91000FF",
      x"FB402702",
      x"C6622500",
      x"30605741",
      x"0203BFFF",
      x"02A41A03",
      x"0B029E07",
      x"3F0204CF",
      x"FF0BEA1A",
      x"01B36CFF",
      x"1000705C",
      x"30AA59F0",
      x"FF70010B",
      x"E91D00D4",
      x"C8FA0F02",
      x"6300B601",
      x"DB00FC40",
      x"540000FE",
      x"609B0260",
      x"305C8D02",
      x"B107DF5F",
      x"20028F00",
      x"00B601D3",
      x"03309FFF",
      x"E08BC1F5",
      x"02CB4203",
      x"DA02DFD5",
      x"2A9A00BF",
      x"9601C4BF",
      x"209A0190",
      x"AB1A9E11",
      x"007D9A00",
      x"2903BF9E",
      x"000C00EF",
      x"FE00006E",
      x"FB0001BF",
      x"003C09EF",
      x"917B00D7",
      x"9103F08B",
      x"0021109F",
      x"DBA74000",
      x"FFFDB700",
      x"FFFD9008",
      x"1B64009E",
      x"FF20FFFA",
      x"22F95009",
      x"FE000122",
      x"15ABDE10",
      x"129C5E03",
      x"EF4CFFD9",
      x"00FF7A01",
      x"3E702001",
      x"00352222",
      x"00EF02B0",
      x"07002A03",
      x"600B008D",
      x"500F10BF",
      x"4410013F",
      x"B80A1BFF",
      x"039CFFFE",
      x"A403CDA1",
      x"FB9902BE",
      x"A2002CFF",
      x"00135951",
      x"BF210000",
      x"FFFA003A",
      x"0003AF2D",
      x"7A000A76",
      x"011D7E10",
      x"7F608553",
      x"3AFFFF51",
      x"11AA9A01",
      x"03BB580B",
      x"69003466",
      x"00009C40",
      x"8ABB15BA",
      x"3AFA0301",
      x"01EC7F13",
      x"04B758C8",
      x"0B044007",
      x"4453B931",
      x"CB920B00",
      x"380350BC",
      x"031F04B5",
      x"BFFF003F",
      x"4BFFDA99",
      x"FD408000",
      x"004BD951",
      x"08DF2220",
      x"F500D06A",
      x"009F0300",
      x"0B00AF07",
      x"70D040BF",
      x"A81002BF",
      x"C0B66FFF",
      x"3D011B00",
      x"FFDBBDFF",
      x"844837DF",
      x"2000BF41",
      x"ABBB0C02",
      x"4B049505",
      x"A701119D",
      x"CB820497",
      x"01A08714",
      x"AA32AE3F",
      x"BA400345",
      x"C8AB30CC",
      x"9F449B04",
      x"FEA99AFF",
      x"1002FF0D",
      x"141F64FA",
      x"66024B17",
      x"A31A0280",
      x"FB4005CF",
      x"019007DF",
      x"74D80960",
      x"0112213F",
      x"CEEC10A6",
      x"FF7D10AB",
      x"709229EF",
      x"50E301FF",
      x"989D527F",
      x"B3599999",
      x"10AFFF04",
      x"AFBB0103",
      x"232014D7",
      x"FFF00163",
      x"FFFBBBB2",
      x"F91B05F3",
      x"13500310",
      x"8F125E22",
      x"BBDF9312",
      x"FF3C5301",
      x"500320DF",
      x"137F2313",
      x"0FFFA063",
      x"FFDBBBA0",
      x"0320DE01",
      x"7F131350",
      x"206313DF",
      x"3F20EF03",
      x"1340AA42",
      x"3A437F13",
      x"00EE049C",
      x"A3034007",
      x"00CC044D",
      x"2705ACE9",
      x"A12B05B4",
      x"57222F05",
      x"002AFFFE",
      x"08033040",
      x"030A7A03",
      x"03AB2B7E",
      x"86036D82",
      x"9E8A039D",
      x"03202731",
      x"336753DD",
      x"CF01506F",
      x"87137F13",
      x"7F3B1200",
      x"236753E9",
      x"2077136F",
      x"03F303EB",
      x"68F7331F",
      x"8003F0BF",
      x"6305A107",
      x"44EFFC30",
      x"4B830508",
      x"CF01B200",
      x"DF69FD50",
      x"77065A00",
      x"707B06B3",
      x"564B03FF",
      x"7C4F034C",
      x"109C5303",
      x"9C7F0603",
      x"7C8206A8",
      x"064C8606",
      x"FFFC1C8A",
      x"FD08EF17",
      x"00FE0300",
      x"20960607",
      x"0F10EF07",
      x"C7051710",
      x"04E73009",
      x"0103E0A3",
      x"3E04A503",
      x"EF7202EF",
      x"BAD406B9",
      x"10B00370",
      x"A004EF0F",
      x"0BFF5F13",
      x"00B15000",
      x"03F00003",
      x"99990B30",
      x"FD431319",
      x"0B4003F0",
      x"03076B03",
      x"0B5003F0",
      x"DF431310",
      x"0B6003F0",
      x"05F30408",
      x"4003F065",
      x"DD43130B",
      x"078003F0",
      x"F083076F",
      x"F90B6003",
      x"F8715F01",
      x"03F0E500",
      x"00000B30",
      x"590308F5",
      x"F10708F2",
      x"0F0003F0",
      x"C50419FF",
      x"F104496A",
      x"08691913",
      x"2408691C",
      x"2508B749",
      x"027D1129",
      x"03087F78",
      x"0B3003F0",
      x"D6A305BF",
      x"03F06407",
      x"4B930770",
      x"5F8303F0",
      x"A303F0FF",
      x"C303F05F",
      x"3603F05F",
      x"062743DF",
      x"00FF1C72",
      x"15370380",
      x"00280897",
      x"5733FAC5",
      x"2F132753",
      x"27183713",
      x"1BCE065D",
      x"065743DA",
      x"E413C4D9",
      x"D6206F48",
      x"FF25FFE9",
      x"AF23096D",
      x"076F0800",
      x"04A47718",
      x"A603AE53",
      x"440640FF",
      x"F8D9D800",
      x"191717DF",
      x"2007A713",
      x"DFF64AFF",
      x"B0B817E3",
      x"4473B35F",
      x"6CD73444",
      x"17B60316",
      x"9FF090B7",
      x"100CBF29",
      x"0CFA0903",
      x"0C170986",
      x"A8444443",
      x"1B030596",
      x"FFFEA100",
      x"FEC9209E",
      x"60000BEF",
      x"6606DCBA",
      x"04CDA733",
      x"CF068073",
      x"DFFEDDDF",
      x"0DBDFF4A",
      x"2344017A",
      x"EF77D917",
      x"63D3064C",
      x"26D74607",
      x"444430DF",
      x"73C33FA8",
      x"607DB0EC",
      x"427B93BF",
      x"73B35FB1",
      x"CADD4444",
      x"4473D3F2",
      x"73D37FB0",
      x"B843A908",
      x"73B38CDF",
      x"B0303444",
      x"4473C3BF",
      x"EBB8DA14",
      x"C14173D3",
      x"4073F35F",
      x"80091FB1",
      x"90094909",
      x"1009FFFE",
      x"4D089CC9",
      x"5EB14460",
      x"3B0BE309",
      x"710429EF",
      x"EDDEFFFF",
      x"21BDAB0B",
      x"A1444335",
      x"AFFF039F",
      x"0BAFAF08",
      x"0AAF41D6",
      x"4442AFF7",
      x"8DB92444",
      x"C073D3FB",
      x"F273C37F",
      x"2073D35E",
      x"73C3DFB1",
      x"C0D04470",
      x"A71201F0",
      x"710000C7",
      x"2000FC03",
      x"0B10FFD9",
      x"AA471AAC",
      x"0AAEDE06",
      x"A20C5C57",
      x"03670A0A",
      x"2A2B08FD",
      x"F2131777",
      x"079F9232",
      x"E71C100B",
      x"EB1CA264",
      x"8100F70C",
      x"16BEBFAA",
      x"ADC30C96",
      x"ACF60C16",
      x"FF1CFA1C",
      x"040DC6A4",
      x"20000F1D",
      x"30EF02A7",
      x"00872852",
      x"AAABEF59",
      x"DDEDDC89",
      x"8C1FF08F",
      x"A8A61F6A",
      x"ADD51CAA",
      x"BA00EF2F",
      x"0AA46C00",
      x"1D194050",
      x"DC09AD77",
      x"BFFF0307",
      x"39BD0039",
      x"F30AC31B",
      x"BFD808B4",
      x"A60C8A0B",
      x"00D0FD00",
      x"12F0D394",
      x"09BA0770",
      x"7D4431CC",
      x"C0FFF38F",
      x"1FE0AFBD",
      x"559ABDEF",
      x"F1D83445",
      x"160A40B4",
      x"01A012F0",
      x"01920000",
      x"04B50323",
      x"07D50645",
      x"0AF10964",
      x"0E050C7C",
      x"11110F8C",
      x"14131294",
      x"1708158F",
      x"19EF187D",
      x"1CC61B5D",
      x"1F8B1E2B",
      x"223D20E7",
      x"24DA238E",
      x"275F261F",
      x"29CD2899",
      x"2C212AFA",
      x"2E5A2D41",
      x"30762F6B",
      x"32743179",
      x"34533367",
      x"36123536",
      x"37AF36E5",
      x"392A3871",
      x"3A8239DA",
      x"3BB63B20",
      x"3CC53C42",
      x"3DAE3D3E",
      x"3E713E14",
      x"3F0E3EC5",
      x"3F843F4E",
      x"3FD33FB1",
      x"3FFB3FEC",
      x"3FFB4000",
      x"3FD33FEC",
      x"3F843FB1",
      x"3F0E3F4E",
      x"3E713EC5",
      x"3DAE3E14",
      x"3CC53D3E",
      x"3BB63C42",
      x"3A823B20",
      x"392A39DA",
      x"37AF3871",
      x"361236E5",
      x"34533536",
      x"32743367",
      x"30763179",
      x"2E5A2F6B",
      x"2C212D41",
      x"29CD2AFA",
      x"275F2899",
      x"24DA261F",
      x"223D238E",
      x"1F8B20E7",
      x"1CC61E2B",
      x"19EF1B5D",
      x"1708187D",
      x"1413158F",
      x"11111294",
      x"0E050F8C",
      x"0AF10C7C",
      x"07D50964",
      x"04B50645",
      x"01920323",
      x"FE6E0000",
      x"FB4BFCDD",
      x"F82BF9BB",
      x"F50FF69C",
      x"F1FBF384",
      x"EEEFF074",
      x"EBEDED6C",
      x"E8F8EA71",
      x"E611E783",
      x"E33AE4A3",
      x"E075E1D5",
      x"DDC3DF19",
      x"DB26DC72",
      x"D8A1D9E1",
      x"D633D767",
      x"D3DFD506",
      x"D1A6D2BF",
      x"CF8AD095",
      x"CD8CCE87",
      x"CBADCC99",
      x"C9EECACA",
      x"C851C91B",
      x"C6D6C78F",
      x"C57EC626",
      x"C44AC4E0",
      x"C33BC3BE",
      x"C252C2C2",
      x"C18FC1EC",
      x"C0F2C13B",
      x"C07CC0B2",
      x"C02DC04F",
      x"C005C014",
      x"C005C000",
      x"C02DC014",
      x"C07CC04F",
      x"C0F2C0B2",
      x"C18FC13B",
      x"C252C1EC",
      x"C33BC2C2",
      x"C44AC3BE",
      x"C57EC4E0",
      x"C6D6C626",
      x"C851C78F",
      x"C9EEC91B",
      x"CBADCACA",
      x"CD8CCC99",
      x"CF8ACE87",
      x"D1A6D095",
      x"D3DFD2BF",
      x"D633D506",
      x"D8A1D767",
      x"DB26D9E1",
      x"DDC3DC72",
      x"E075DF19",
      x"E33AE1D5",
      x"E611E4A3",
      x"E8F8E783",
      x"EBEDEA71",
      x"EEEFED6C",
      x"F1FBF074",
      x"F50FF384",
      x"F82BF69C",
      x"FB4BF9BB",
      x"FE6EFCDD",
      x"E3E2E1E0",
      x"E7E6E5E4",
      x"EBEAE9E8",
      x"D3D2D1D0",
      x"D7D6D5D4",
      x"DBDAD9D8",
      x"C3C2C1C0",
      x"C7C6C5C4",
      x"CBCAC9C8",
      x"B3B2B1B0",
      x"B7B6B5B4",
      x"BBBAB9B8",
      x"A3A2A1A0",
      x"A7A6A5A4",
      x"ABAAA9A8",
      x"93929190",
      x"97969594",
      x"9B9A9998",
      x"83828180",
      x"87868584",
      x"8B8A8988",
      x"73727170",
      x"77767574",
      x"7B7A7978",
      x"63626160",
      x"67666564",
      x"6B6A6968",
      x"53525150",
      x"57565554",
      x"5B5A5958",
      x"43424140",
      x"47464544",
      x"4B4A4948",
      x"33323130",
      x"37363534",
      x"3B3A3938",
      x"23222120",
      x"27262524",
      x"2B2A2928",
      x"13121110",
      x"17161514",
      x"1B1A1918",
      x"03020100",
      x"07060504",
      x"0B0A0908",
      x"80000000",
      x"879C7C97",
      x"8FACD61E",
      x"9837F052",
      x"A14517CC",
      x"AADC0848",
      x"B504F334",
      x"BFC886BB",
      x"CB2FF52A",
      x"D744FCCB",
      x"E411F03A",
      x"F1A1BF39",
      x"52416B64",
      x"0000004D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(to_integer(unsigned(address)));
      end if;
   end process;

   process (clk) 
   begin
      if rising_edge(clk) then
         if wren = '1' then
            rom(to_integer(unsigned(wraddress))) <= wrdata;
         end if;
      end if;
   end process;

end architecture;
